Require Export premises.

Set Implicit Arguments.
Unset Strict Implicit.
Unset Printing Implicit Defensive.

(** The module to deal with finite or infinite sequences. *)
Module Sequence.



End Sequence.